`timescale 1ps/1ps

module hazardunit(
    clk,
    RegWriteW, 
    RegWriteM,  
    ForwardAE, 
    ForwardBE,
    Match_1E_M,
    Match_1E_W,
    Match_2E_M,
    Match_2E_W
);






endmodule