`timescale 1ns / 1ps

module basysdecoder (
    output reg [6:0] out0,        
    output wire [3:0] enable,      
    input wire clk,               
    input wire real_clk,         
    input wire [15:0] ResultW 
);

    reg [1:0] state;             
    reg [3:0] digito;            
    reg activo;                 

    assign enable = 4'b0000;

    localparam S0 = 2'b00;       
    localparam S1 = 2'b01;       
    localparam S2 = 2'b10;       
    localparam S3 = 2'b11;       

    always @(posedge clk or posedge real_clk) begin
        if (real_clk)
        begin
            state <= S0;
            activo <= 1;
        end
        else if (activo) 
        begin
            case (state)
                S0: state <= S1;
                S1: state <= S2;
                S2: state <= S3;
                S3: activo <= 0; 
            endcase
        end 
         
    end

    always @(*) begin
        case (state)
            S0: digito = ResultW[3:0];    
            S1: digito = ResultW[7:4];    
            S2: digito = ResultW[11:8];   
            S3: digito = ResultW[15:12];  
            default: digito = 4'b0000;
        endcase
    end

    always @(*) begin
        case (digito)
            4'b0000: out0 = 7'b0000001; // 0
            4'b0001: out0 = 7'b1001111; // 1
            4'b0010: out0 = 7'b0010010; // 2
            4'b0011: out0 = 7'b0000110; // 3
            4'b0100: out0 = 7'b1001100; // 4
            4'b0101: out0 = 7'b0100100; // 5
            4'b0110: out0 = 7'b0100000; // 6
            4'b0111: out0 = 7'b0001111; // 7
            4'b1000: out0 = 7'b0000000; // 8
            4'b1001: out0 = 7'b0001100; // 9
            4'b1010: out0 = 7'b0001000; // A
            4'b1011: out0 = 7'b1100000; // b
            4'b1100: out0 = 7'b0110001; // C
            4'b1101: out0 = 7'b1000010; // d
            4'b1110: out0 = 7'b0110000; // E
            4'b1111: out0 = 7'b0111000; // F
            default: out0 = 7'b1111111; // Default (all segments off)
        endcase
    end

endmodule
